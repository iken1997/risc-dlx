LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY FA IS
  PORT (
    A : IN STD_LOGIC;
    B : IN STD_LOGIC;
    Ci : IN STD_LOGIC;
    S : OUT STD_LOGIC;
    Co : OUT STD_LOGIC);
END FA;

ARCHITECTURE BEHAVIORAL OF FA IS

BEGIN

  S <= A XOR B XOR Ci;
  Co <= (A AND B) OR (B AND Ci) OR (A AND Ci);

END BEHAVIORAL;
