LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.std_logic_arith.ALL;
USE work.CONSTANTS.ALL;

ENTITY DLX_TestBench IS
	GENERIC (
		FILENAME : STRING := "Branch.mem"--"test-arith.mem" -- change filename to change asm test
	);
END DLX_TestBench;

ARCHITECTURE tb OF DLX_TestBench IS

	COMPONENT IRAM IS
		GENERIC (
			FILENAME  : STRING  := "test.asm.mem";
			RAM_DEPTH : INTEGER := 128;
			I_SIZE    : INTEGER := 32);
		PORT (
			Rst  : IN STD_LOGIC;
			EN   : STD_LOGIC;
			RDY  : STD_LOGIC;
			Addr : IN STD_LOGIC_VECTOR(I_SIZE - 1 DOWNTO 0);
			Dout : OUT STD_LOGIC_VECTOR(I_SIZE - 1 DOWNTO 0)
		);

	END COMPONENT;

	COMPONENT DRAM IS
		GENERIC (
			MEM_SIZE : INTEGER := 512;
			NADD     : INTEGER := 6
		);
		PORT (
			DATA_IN  : IN WORD;
			DATA_OUT : OUT WORD;
			ADDR     : IN STD_LOGIC_VECTOR (NADD - 1 DOWNTO 0);
			EN       : STD_LOGIC;
			RDY      : STD_LOGIC;
			R_EN     : STD_LOGIC;
			W_EN     : STD_LOGIC;
			CLK      : STD_LOGIC;
			RST      : STD_LOGIC
		);
	END COMPONENT;

	COMPONENT DLX IS
		GENERIC (
			IR_SIZE : INTEGER := 32; -- Instruction Register Size
			PC_SIZE : INTEGER := 32  -- Program Counter Size
		);
		PORT (
			-- Inputs
			CLK : IN STD_LOGIC; -- Clock
			RST : IN STD_LOGIC; -- Reset:Active-High

			IRAM_ADDRESS : OUT STD_LOGIC_VECTOR(IR_SIZE - 1 DOWNTO 0);
			IRAM_ISSUE   : OUT STD_LOGIC;
			IRAM_READY   : IN STD_LOGIC;
			IRAM_DATA    : IN STD_LOGIC_VECTOR (WORD_SIZE - 1 DOWNTO 0);

			DRAM_ADDRESS  : OUT STD_LOGIC_VECTOR(IR_SIZE - 1 DOWNTO 0);
			DRAM_ISSUE    : OUT STD_LOGIC;
			DRAM_READ     : OUT STD_LOGIC;
			DRAM_WRITE    : OUT STD_LOGIC;
			DRAM_READY    : IN STD_LOGIC;
			DRAM_DATA_OUT : IN STD_LOGIC_VECTOR (WORD_SIZE - 1 DOWNTO 0);
			DRAM_DATA_IN  : OUT STD_LOGIC_VECTOR (WORD_SIZE - 1 DOWNTO 0)
		);
	END COMPONENT;

	SIGNAL CLK          : STD_LOGIC := '0'; -- Clock
	SIGNAL RST          : STD_LOGIC;        -- Reset:Active-Low
	SIGNAL IRAM_ADDRESS : STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);
	SIGNAL PC           : STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);
	SIGNAL IRAM_ENABLE  : STD_LOGIC;
	SIGNAL IRAM_READY   : STD_LOGIC;
	SIGNAL IRAM_DATA    : STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);

	SIGNAL DRAM_ADDRESS  : STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);
	SIGNAL DRAM_ENABLE   : STD_LOGIC;
	SIGNAL DRAM_READ     : STD_LOGIC;
	SIGNAL DRAM_WRITE    : STD_LOGIC;
	SIGNAL DRAM_READY    : STD_LOGIC;
	SIGNAL DRAM_DATA_IN  : STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);
	SIGNAL DRAM_DATA_OUT : STD_LOGIC_VECTOR(WORD_SIZE - 1 DOWNTO 0);

BEGIN
  IRAM_ADDRESS <=  "00" & PC(PC'left DOWNTO PC'right +2); 
	-- IRAM
	INSTR_RAM : IRAM
	GENERIC MAP(
		FILENAME  => FILENAME,
		RAM_DEPTH => 128,
		I_SIZE    => 32
	)
	PORT MAP(
		Rst  => Rst,
		EN   => IRAM_ENABLE,
		RDY  => IRAM_READY,
		Addr => IRAM_ADDRESS,
		Dout => IRAM_DATA
	);
	-- DRAM
	DATA_RAM : DRAM
	GENERIC MAP(
		MEM_SIZE => DRAM_SIZE,
		NADD     => WORD_SIZE
	)
	PORT MAP(
		DATA_IN  => DRAM_DATA_IN,
		DATA_OUT => DRAM_DATA_OUT,
		ADDR     => DRAM_ADDRESS,
		EN       => DRAM_ENABLE,
		RDY      => DRAM_READY,
		R_EN     => DRAM_READ,
		W_EN     => DRAM_WRITE,
		CLK      => CLK,
		RST      => RST
	);

	-- DLX
	dlx_inst : DLX
	GENERIC MAP(
		IR_SIZE => WORD_SIZE,
		PC_SIZE => WORD_SIZE
	)
	PORT MAP(
		CLK           => CLK,
		RST           => RST,
		IRAM_ADDRESS  => PC,
		IRAM_ISSUE    => IRAM_ENABLE,
		IRAM_READY    => IRAM_READY,
		IRAM_DATA     => IRAM_DATA,
		DRAM_ADDRESS  => DRAM_ADDRESS,
		DRAM_ISSUE    => DRAM_ENABLE,
		DRAM_READ     => DRAM_READ,
		DRAM_WRITE    => DRAM_WRITE,
		DRAM_READY    => DRAM_READY,
		DRAM_DATA_OUT => DRAM_DATA_OUT,
		DRAM_DATA_IN  => DRAM_DATA_IN
	);

	Clk <= NOT Clk AFTER 10 ns;
	Rst <= '0', '1' AFTER 12 ns;

END tb;
