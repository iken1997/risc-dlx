LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;
USE ieee.math_real.ALL;
USE ieee.std_logic_unsigned.ALL;
USE ieee.std_logic_arith.ALL;
USE WORK.myTypes.ALL;
USE WORK.CONSTANTS.ALL;
PACKAGE alu_types IS
	TYPE TYPE_OP IS (NOP, ADD, SUB, MULT, BITAND, BITOR, BITXOR, BITNOT, FUNCLSL, FUNCLSR, FUNCRL, FUNCRR, GREATER_EQ, UGREATER_EQ, LOWER_EQ, ULOWER_EQ, EQ, NEQ);

	FUNCTION func_decode (vector : STD_LOGIC_VECTOR) RETURN TYPE_OP;

END alu_types;

PACKAGE BODY alu_types IS

	FUNCTION func_decode (vector : STD_LOGIC_VECTOR) RETURN TYPE_OP IS
		VARIABLE FUNC : TYPE_OP;
	BEGIN
		CASE conv_integer(vector) IS
			WHEN 0 => FUNC := NOP;
			WHEN 1 => FUNC := ADD;
			WHEN 2 => FUNC := SUB;
			WHEN 3 => FUNC := MULT;
			WHEN 4 => FUNC := BITAND;
			WHEN 5 => FUNC := BITOR;
			WHEN 6 => FUNC := BITXOR;
			WHEN 7 => FUNC := BITNOT;
			WHEN 8 => FUNC := FUNCLSL;
			WHEN 9 => FUNC := FUNCLSR;
			WHEN 10 => FUNC := FUNCRL;
			WHEN 11 => FUNC := FUNCRR;
			WHEN 12 => FUNC := GREATER_EQ;
			WHEN 13 => FUNC := UGREATER_EQ;
			WHEN 14 => FUNC := LOWER_EQ;
			WHEN 15 => FUNC := ULOWER_EQ;
			WHEN 16 => FUNC := EQ;
			WHEN 17 => FUNC := NEQ;
			WHEN OTHERS => FUNC := NOP;
		END CASE;
		RETURN FUNC;
	END FUNCTION func_decode;

END PACKAGE BODY alu_types;
