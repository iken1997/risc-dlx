LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE WORK.CONSTANTS.all;

ENTITY MUX21_GENERIC IS
GENERIC (
	NBIT : INTEGER := NumBit);
PORT (
	A : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
	B : IN STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0);
	SEL : IN STD_LOGIC;
	Y : OUT STD_LOGIC_VECTOR(NBIT - 1 DOWNTO 0));
END MUX21_GENERIC;
ARCHITECTURE behavioral OF MUX21_GENERIC IS
BEGIN
WITH SEL SELECT
	Y <= A WHEN '0',
	B WHEN OTHERS;
END behavioral;

ARCHITECTURE structural OF MUX21_GENERIC IS
COMPONENT MUX21
	PORT (
		A : IN STD_LOGIC;
		B : IN STD_LOGIC;
		SEL : IN STD_LOGIC;
		Y : OUT STD_LOGIC);
END COMPONENT;
BEGIN
g1 : FOR i IN 0 TO NBIT - 1 GENERATE
	MUX : MUX21 PORT MAP(A => A(i), B => B(i), SEL => SEL, Y => Y(i));
END GENERATE;
END structural;

CONFIGURATION CFG_MUX21_GEN_BEHAVIORAL OF MUX21_GENERIC IS
FOR BEHAVIORAL
END FOR;
END CFG_MUX21_GEN_BEHAVIORAL;

CONFIGURATION CFG_MUX21_GEN_STRUCTURAL OF MUX21_GENERIC IS
FOR STRUCTURAL
END FOR;
END CFG_MUX21_GEN_STRUCTURAL;